// Test file for IP-XACT conversion
// See test_samples/LICENSE.md for license information


module test_various_patterns (
    input  wire        clk,
    input  wire        rst_n,

    // Pattern 1: Standard M_AXI_AWADDR
    output wire [31:0] M_AXI_AWADDR,
    output wire [7:0]  M_AXI_AWLEN,
    output wire [2:0]  M_AXI_AWSIZE,
    output wire [1:0]  M_AXI_AWBURST,
    output wire        M_AXI_AWVALID,
    input  wire        M_AXI_AWREADY,
    output wire [31:0] M_AXI_WDATA,
    output wire [3:0]  M_AXI_WSTRB,
    output wire        M_AXI_WLAST,
    output wire        M_AXI_WVALID,
    input  wire        M_AXI_WREADY,
    input  wire [1:0]  M_AXI_BRESP,
    input  wire        M_AXI_BVALID,
    output wire        M_AXI_BREADY,
    output wire [31:0] M_AXI_ARADDR,
    output wire [7:0]  M_AXI_ARLEN,
    output wire [2:0]  M_AXI_ARSIZE,
    output wire [1:0]  M_AXI_ARBURST,
    output wire        M_AXI_ARVALID,
    input  wire        M_AXI_ARREADY,
    input  wire [31:0] M_AXI_RDATA,
    input  wire [1:0]  M_AXI_RRESP,
    input  wire        M_AXI_RLAST,
    input  wire        M_AXI_RVALID,
    output wire        M_AXI_RREADY,

    // Pattern 2: With postfix _o and _i
    output wire [31:0] M_AXI_AWADDR_o,
    output wire [7:0]  M_AXI_AWLEN_o,
    output wire [2:0]  M_AXI_AWSIZE_o,
    output wire [1:0]  M_AXI_AWBURST_o,
    output wire        M_AXI_AWVALID_o,
    input  wire        M_AXI_AWREADY_i,
    output wire [31:0] M_AXI_WDATA_o,
    output wire [3:0]  M_AXI_WSTRB_o,
    output wire        M_AXI_WLAST_o,
    output wire        M_AXI_WVALID_o,
    input  wire        M_AXI_WREADY_i,
    input  wire [1:0]  M_AXI_BRESP_i,
    input  wire        M_AXI_BVALID_i,
    output wire        M_AXI_BREADY_o,
    output wire [31:0] M_AXI_ARADDR_o,
    output wire [7:0]  M_AXI_ARLEN_o,
    output wire [2:0]  M_AXI_ARSIZE_o,
    output wire [1:0]  M_AXI_ARBURST_o,
    output wire        M_AXI_ARVALID_o,
    input  wire        M_AXI_ARREADY_i,
    input  wire [31:0] M_AXI_RDATA_i,
    input  wire [1:0]  M_AXI_RRESP_i,
    input  wire        M_AXI_RLAST_i,
    input  wire        M_AXI_RVALID_i,
    output wire        M_AXI_RREADY_o,

    // Pattern 3: Lowercase prefix m_axi_awaddr
    output wire [31:0] m_axi_awaddr,
    output wire [7:0]  m_axi_awlen,
    output wire [2:0]  m_axi_awsize,
    output wire [1:0]  m_axi_awburst,
    output wire        m_axi_awvalid,
    input  wire        m_axi_awready,
    output wire [31:0] m_axi_wdata,
    output wire [3:0]  m_axi_wstrb,
    output wire        m_axi_wlast,
    output wire        m_axi_wvalid,
    input  wire        m_axi_wready,
    input  wire [1:0]  m_axi_bresp,
    input  wire        m_axi_bvalid,
    output wire        m_axi_bready,
    output wire [31:0] m_axi_araddr,
    output wire [7:0]  m_axi_arlen,
    output wire [2:0]  m_axi_arsize,
    output wire [1:0]  m_axi_arburst,
    output wire        m_axi_arvalid,
    input  wire        m_axi_arready,
    input  wire [31:0] m_axi_rdata,
    input  wire [1:0]  m_axi_rresp,
    input  wire        m_axi_rlast,
    input  wire        m_axi_rvalid,
    output wire        m_axi_rready,

    // Pattern 4: With instance number M_AXI0_AWADDR
    output wire [31:0] M_AXI0_AWADDR,
    output wire [7:0]  M_AXI0_AWLEN,
    output wire [2:0]  M_AXI0_AWSIZE,
    output wire [1:0]  M_AXI0_AWBURST,
    output wire        M_AXI0_AWVALID,
    input  wire        M_AXI0_AWREADY,
    output wire [31:0] M_AXI0_WDATA,
    output wire [3:0]  M_AXI0_WSTRB,
    output wire        M_AXI0_WLAST,
    output wire        M_AXI0_WVALID,
    input  wire        M_AXI0_WREADY,
    input  wire [1:0]  M_AXI0_BRESP,
    input  wire        M_AXI0_BVALID,
    output wire        M_AXI0_BREADY,
    output wire [31:0] M_AXI0_ARADDR,
    output wire [7:0]  M_AXI0_ARLEN,
    output wire [2:0]  M_AXI0_ARSIZE,
    output wire [1:0]  M_AXI0_ARBURST,
    output wire        M_AXI0_ARVALID,
    input  wire        M_AXI0_ARREADY,
    input  wire [31:0] M_AXI0_RDATA,
    input  wire [1:0]  M_AXI0_RRESP,
    input  wire        M_AXI0_RLAST,
    input  wire        M_AXI0_RVALID,
    output wire        M_AXI0_RREADY
);

endmodule
